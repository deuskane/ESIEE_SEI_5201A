library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std   .all;

entity labo01 is
  
end entity labo01;

architecture rtl of labo01 is

begin  -- architecture rtl

end architecture rtl;
